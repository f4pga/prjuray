// Copyright 2020-2022 F4PGA Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// SPDX-License-Identifier: Apache-2.0

module top(input clk, stb, di, output do);
	roi roi(
		.clk(clk),
		.stb(stb),
		.di(di),
		.do(do)
	);
endmodule

module roi(input clk, stb, di, output do);
	reg do_reg = 0;
	always @(posedge clk) begin
		if (stb) begin
			do_reg <= di;
		end
	end
	assign do = do_reg;
endmodule
