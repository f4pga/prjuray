module top(
    output wire [1:0] led
);

    wire pl_clk3,pl_clk2,pl_clk1,pl_clk_unbuffered;

    localparam BITS = 2;
    localparam LOG2DELAY = 24;

    reg [BITS+LOG2DELAY-1:0] counter = 0;

    always @(posedge pl_clk0) begin
        counter <= counter + 1;
    end

    assign led = counter >> LOG2DELAY;

  (* BOX_TYPE = "PRIMITIVE" *)
  (* KEEP, DONT_TOUCH *)
  PS8 PS8_i
       (.ADMA2PLCACK(),
        .ADMA2PLTVLD(),
        .ADMAFCICLK(),
        .AIBPMUAFIFMFPDACK(),
        .AIBPMUAFIFMLPDACK(),
        .DDRCEXTREFRESHRANK0REQ(),
        .DDRCEXTREFRESHRANK1REQ(),
        .DDRCREFRESHPLCLK(),
        .DPAUDIOREFCLK(),
        .DPAUXDATAIN(),
        .DPAUXDATAOEN(),
        .DPAUXDATAOUT(),
        .DPEXTERNALCUSTOMEVENT1(),
        .DPEXTERNALCUSTOMEVENT2(),
        .DPEXTERNALVSYNCEVENT(),
        .DPHOTPLUGDETECT(),
        .DPLIVEGFXALPHAIN(),
        .DPLIVEGFXPIXEL1IN(),
        .DPLIVEVIDEODEOUT(),
        .DPLIVEVIDEOINDE(),
        .DPLIVEVIDEOINHSYNC(),
        .DPLIVEVIDEOINPIXEL1(),
        .DPLIVEVIDEOINVSYNC(),
        .DPMAXISMIXEDAUDIOTDATA(),
        .DPMAXISMIXEDAUDIOTID(),
        .DPMAXISMIXEDAUDIOTREADY(),
        .DPMAXISMIXEDAUDIOTVALID(),
        .DPSAXISAUDIOCLK(),
        .DPSAXISAUDIOTDATA(),
        .DPSAXISAUDIOTID(),
        .DPSAXISAUDIOTREADY(),
        .DPSAXISAUDIOTVALID(),
        .DPVIDEOINCLK(),
        .DPVIDEOOUTHSYNC(),
        .DPVIDEOOUTPIXEL1(),
        .DPVIDEOOUTVSYNC(),
        .DPVIDEOREFCLK(),
        .EMIOCAN0PHYRX(),
        .EMIOCAN0PHYTX(),
        .EMIOCAN1PHYRX(),
        .EMIOCAN1PHYTX(),
        .EMIOENET0DMABUSWIDTH(),
        .EMIOENET0DMATXENDTOG(),
        .EMIOENET0DMATXSTATUSTOG(),
        .EMIOENET0EXTINTIN(),
        .EMIOENET0GEMTSUTIMERCNT(),
        .EMIOENET0GMIICOL(),
        .EMIOENET0GMIICRS(),
        .EMIOENET0GMIIRXCLK(),
        .EMIOENET0GMIIRXD(),
        .EMIOENET0GMIIRXDV(),
        .EMIOENET0GMIIRXER(),
        .EMIOENET0GMIITXCLK(),
        .EMIOENET0GMIITXD(),
        .EMIOENET0GMIITXEN(),
        .EMIOENET0GMIITXER(),
        .EMIOENET0MDIOI(),
        .EMIOENET0MDIOMDC(),
        .EMIOENET0MDIOO(),
        .EMIOENET0MDIOTN(),
        .EMIOENET0RXWDATA(),
        .EMIOENET0RXWEOP(),
        .EMIOENET0RXWERR(),
        .EMIOENET0RXWFLUSH(),
        .EMIOENET0RXWOVERFLOW(),
        .EMIOENET0RXWSOP(),
        .EMIOENET0RXWSTATUS(),
        .EMIOENET0RXWWR(),
        .EMIOENET0SPEEDMODE(),
        .EMIOENET0TXRCONTROL(),
        .EMIOENET0TXRDATA(),
        .EMIOENET0TXRDATARDY(),
        .EMIOENET0TXREOP(),
        .EMIOENET0TXRERR(),
        .EMIOENET0TXRFLUSHED(),
        .EMIOENET0TXRRD(),
        .EMIOENET0TXRSOP(),
        .EMIOENET0TXRSTATUS(),
        .EMIOENET0TXRUNDERFLOW(),
        .EMIOENET0TXRVALID(),
        .EMIOENET1DMABUSWIDTH(),
        .EMIOENET1DMATXENDTOG(),
        .EMIOENET1DMATXSTATUSTOG(),
        .EMIOENET1EXTINTIN(),
        .EMIOENET1GMIICOL(),
        .EMIOENET1GMIICRS(),
        .EMIOENET1GMIIRXCLK(),
        .EMIOENET1GMIIRXD(),
        .EMIOENET1GMIIRXDV(),
        .EMIOENET1GMIIRXER(),
        .EMIOENET1GMIITXCLK(),
        .EMIOENET1GMIITXD(),
        .EMIOENET1GMIITXEN(),
        .EMIOENET1GMIITXER(),
        .EMIOENET1MDIOI(),
        .EMIOENET1MDIOMDC(),
        .EMIOENET1MDIOO(),
        .EMIOENET1MDIOTN(),
        .EMIOENET1RXWDATA(),
        .EMIOENET1RXWEOP(),
        .EMIOENET1RXWERR(),
        .EMIOENET1RXWFLUSH(),
        .EMIOENET1RXWOVERFLOW(),
        .EMIOENET1RXWSOP(),
        .EMIOENET1RXWSTATUS(),
        .EMIOENET1RXWWR(),
        .EMIOENET1SPEEDMODE(),
        .EMIOENET1TXRCONTROL(),
        .EMIOENET1TXRDATA(),
        .EMIOENET1TXRDATARDY(),
        .EMIOENET1TXREOP(),
        .EMIOENET1TXRERR(),
        .EMIOENET1TXRFLUSHED(),
        .EMIOENET1TXRRD(),
        .EMIOENET1TXRSOP(),
        .EMIOENET1TXRSTATUS(),
        .EMIOENET1TXRUNDERFLOW(),
        .EMIOENET1TXRVALID(),
        .EMIOENET2DMABUSWIDTH(),
        .EMIOENET2DMATXENDTOG(),
        .EMIOENET2DMATXSTATUSTOG(),
        .EMIOENET2EXTINTIN(),
        .EMIOENET2GMIICOL(),
        .EMIOENET2GMIICRS(),
        .EMIOENET2GMIIRXCLK(),
        .EMIOENET2GMIIRXD(),
        .EMIOENET2GMIIRXDV(),
        .EMIOENET2GMIIRXER(),
        .EMIOENET2GMIITXCLK(),
        .EMIOENET2GMIITXD(),
        .EMIOENET2GMIITXEN(),
        .EMIOENET2GMIITXER(),
        .EMIOENET2MDIOI(),
        .EMIOENET2MDIOMDC(),
        .EMIOENET2MDIOO(),
        .EMIOENET2MDIOTN(),
        .EMIOENET2RXWDATA(),
        .EMIOENET2RXWEOP(),
        .EMIOENET2RXWERR(),
        .EMIOENET2RXWFLUSH(),
        .EMIOENET2RXWOVERFLOW(),
        .EMIOENET2RXWSOP(),
        .EMIOENET2RXWSTATUS(),
        .EMIOENET2RXWWR(),
        .EMIOENET2SPEEDMODE(),
        .EMIOENET2TXRCONTROL(),
        .EMIOENET2TXRDATA(),
        .EMIOENET2TXRDATARDY(),
        .EMIOENET2TXREOP(),
        .EMIOENET2TXRERR(),
        .EMIOENET2TXRFLUSHED(),
        .EMIOENET2TXRRD(),
        .EMIOENET2TXRSOP(),
        .EMIOENET2TXRSTATUS(),
        .EMIOENET2TXRUNDERFLOW(),
        .EMIOENET2TXRVALID(),
        .EMIOENET3DMABUSWIDTH(),
        .EMIOENET3DMATXENDTOG(),
        .EMIOENET3DMATXSTATUSTOG(),
        .EMIOENET3EXTINTIN(),
        .EMIOENET3GMIICOL(),
        .EMIOENET3GMIICRS(),
        .EMIOENET3GMIIRXCLK(),
        .EMIOENET3GMIIRXD(),
        .EMIOENET3GMIIRXDV(),
        .EMIOENET3GMIIRXER(),
        .EMIOENET3GMIITXCLK(),
        .EMIOENET3GMIITXD(),
        .EMIOENET3GMIITXEN(),
        .EMIOENET3GMIITXER(),
        .EMIOENET3MDIOI(),
        .EMIOENET3MDIOMDC(),
        .EMIOENET3MDIOO(),
        .EMIOENET3MDIOTN(),
        .EMIOENET3RXWDATA(),
        .EMIOENET3RXWEOP(),
        .EMIOENET3RXWERR(),
        .EMIOENET3RXWFLUSH(),
        .EMIOENET3RXWOVERFLOW(),
        .EMIOENET3RXWSOP(),
        .EMIOENET3RXWSTATUS(),
        .EMIOENET3RXWWR(),
        .EMIOENET3SPEEDMODE(),
        .EMIOENET3TXRCONTROL(),
        .EMIOENET3TXRDATA(),
        .EMIOENET3TXRDATARDY(),
        .EMIOENET3TXREOP(),
        .EMIOENET3TXRERR(),
        .EMIOENET3TXRFLUSHED(),
        .EMIOENET3TXRRD(),
        .EMIOENET3TXRSOP(),
        .EMIOENET3TXRSTATUS(),
        .EMIOENET3TXRUNDERFLOW(),
        .EMIOENET3TXRVALID(),
        .EMIOENETTSUCLK(),
        .EMIOGEM0DELAYREQRX(),
        .EMIOGEM0DELAYREQTX(),
        .EMIOGEM0PDELAYREQRX(),
        .EMIOGEM0PDELAYREQTX(),
        .EMIOGEM0PDELAYRESPRX(),
        .EMIOGEM0PDELAYRESPTX(),
        .EMIOGEM0RXSOF(),
        .EMIOGEM0SYNCFRAMERX(),
        .EMIOGEM0SYNCFRAMETX(),
        .EMIOGEM0TSUINCCTRL(),
        .EMIOGEM0TSUTIMERCMPVAL(),
        .EMIOGEM0TXRFIXEDLAT(),
        .EMIOGEM0TXSOF(),
        .EMIOGEM1DELAYREQRX(),
        .EMIOGEM1DELAYREQTX(),
        .EMIOGEM1PDELAYREQRX(),
        .EMIOGEM1PDELAYREQTX(),
        .EMIOGEM1PDELAYRESPRX(),
        .EMIOGEM1PDELAYRESPTX(),
        .EMIOGEM1RXSOF(),
        .EMIOGEM1SYNCFRAMERX(),
        .EMIOGEM1SYNCFRAMETX(),
        .EMIOGEM1TSUINCCTRL(),
        .EMIOGEM1TSUTIMERCMPVAL(),
        .EMIOGEM1TXRFIXEDLAT(),
        .EMIOGEM1TXSOF(),
        .EMIOGEM2DELAYREQRX(),
        .EMIOGEM2DELAYREQTX(),
        .EMIOGEM2PDELAYREQRX(),
        .EMIOGEM2PDELAYREQTX(),
        .EMIOGEM2PDELAYRESPRX(),
        .EMIOGEM2PDELAYRESPTX(),
        .EMIOGEM2RXSOF(),
        .EMIOGEM2SYNCFRAMERX(),
        .EMIOGEM2SYNCFRAMETX(),
        .EMIOGEM2TSUINCCTRL(),
        .EMIOGEM2TSUTIMERCMPVAL(),
        .EMIOGEM2TXRFIXEDLAT(),
        .EMIOGEM2TXSOF(),
        .EMIOGEM3DELAYREQRX(),
        .EMIOGEM3DELAYREQTX(),
        .EMIOGEM3PDELAYREQRX(),
        .EMIOGEM3PDELAYREQTX(),
        .EMIOGEM3PDELAYRESPRX(),
        .EMIOGEM3PDELAYRESPTX(),
        .EMIOGEM3RXSOF(),
        .EMIOGEM3SYNCFRAMERX(),
        .EMIOGEM3SYNCFRAMETX(),
        .EMIOGEM3TSUINCCTRL(),
        .EMIOGEM3TSUTIMERCMPVAL(),
        .EMIOGEM3TXRFIXEDLAT(),
        .EMIOGEM3TXSOF(),
        .EMIOGPIOI(),
        .EMIOGPIOO(),
        .EMIOGPIOTN(),
        .EMIOHUBPORTOVERCRNTUSB20(),
        .EMIOHUBPORTOVERCRNTUSB21(),
        .EMIOHUBPORTOVERCRNTUSB30(),
        .EMIOHUBPORTOVERCRNTUSB31(),
        .EMIOI2C0SCLI(),
        .EMIOI2C0SCLO(),
        .EMIOI2C0SCLTN(),
        .EMIOI2C0SDAI(),
        .EMIOI2C0SDAO(),
        .EMIOI2C0SDATN(),
        .EMIOI2C1SCLI(),
        .EMIOI2C1SCLO(),
        .EMIOI2C1SCLTN(),
        .EMIOI2C1SDAI(),
        .EMIOI2C1SDAO(),
        .EMIOI2C1SDATN(),
        .EMIOSDIO0BUSPOWER(),
        .EMIOSDIO0BUSVOLT(),
        .EMIOSDIO0CDN(),
        .EMIOSDIO0CLKOUT(),
        .EMIOSDIO0CMDENA(),
        .EMIOSDIO0CMDIN(),
        .EMIOSDIO0CMDOUT(),
        .EMIOSDIO0DATAENA(),
        .EMIOSDIO0DATAIN(),
        .EMIOSDIO0DATAOUT(),
        .EMIOSDIO0FBCLKIN(),
        .EMIOSDIO0LEDCONTROL(),
        .EMIOSDIO0WP(),
        .EMIOSDIO1BUSPOWER(),
        .EMIOSDIO1BUSVOLT(),
        .EMIOSDIO1CDN(),
        .EMIOSDIO1CLKOUT(),
        .EMIOSDIO1CMDENA(),
        .EMIOSDIO1CMDIN(),
        .EMIOSDIO1CMDOUT(),
        .EMIOSDIO1DATAENA(),
        .EMIOSDIO1DATAIN(),
        .EMIOSDIO1DATAOUT(),
        .EMIOSDIO1FBCLKIN(),
        .EMIOSDIO1LEDCONTROL(),
        .EMIOSDIO1WP(),
        .EMIOSPI0MI(),
        .EMIOSPI0MO(),
        .EMIOSPI0MOTN(),
        .EMIOSPI0SCLKI(),
        .EMIOSPI0SCLKO(),
        .EMIOSPI0SCLKTN(),
        .EMIOSPI0SI(),
        .EMIOSPI0SO(),
        .EMIOSPI0SSIN(),
        .EMIOSPI0SSNTN(),
        .EMIOSPI0SSON(),
        .EMIOSPI0STN(),
        .EMIOSPI1MI(),
        .EMIOSPI1MO(),
        .EMIOSPI1MOTN(),
        .EMIOSPI1SCLKI(),
        .EMIOSPI1SCLKO(),
        .EMIOSPI1SCLKTN(),
        .EMIOSPI1SI(),
        .EMIOSPI1SO(),
        .EMIOSPI1SSIN(),
        .EMIOSPI1SSNTN(),
        .EMIOSPI1SSON(),
        .EMIOSPI1STN(),
        .EMIOTTC0CLKI(),
        .EMIOTTC0WAVEO(),
        .EMIOTTC1CLKI(),
        .EMIOTTC1WAVEO(),
        .EMIOTTC2CLKI(),
        .EMIOTTC2WAVEO(),
        .EMIOTTC3CLKI(),
        .EMIOTTC3WAVEO(),
        .EMIOU2DSPORTVBUSCTRLUSB30(),
        .EMIOU2DSPORTVBUSCTRLUSB31(),
        .EMIOU3DSPORTVBUSCTRLUSB30(),
        .EMIOU3DSPORTVBUSCTRLUSB31(),
        .EMIOUART0CTSN(),
        .EMIOUART0DCDN(),
        .EMIOUART0DSRN(),
        .EMIOUART0DTRN(),
        .EMIOUART0RIN(),
        .EMIOUART0RTSN(),
        .EMIOUART0RX(),
        .EMIOUART0TX(),
        .EMIOUART1CTSN(),
        .EMIOUART1DCDN(),
        .EMIOUART1DSRN(),
        .EMIOUART1DTRN(),
        .EMIOUART1RIN(),
        .EMIOUART1RTSN(),
        .EMIOUART1RX(),
        .EMIOUART1TX(),
        .EMIOWDT0CLKI(),
        .EMIOWDT0RSTO(),
        .EMIOWDT1CLKI(),
        .EMIOWDT1RSTO(),
        .FMIOGEM0FIFORXCLKFROMPL(),
        .FMIOGEM0FIFORXCLKTOPLBUFG(),
        .FMIOGEM0FIFOTXCLKFROMPL(),
        .FMIOGEM0FIFOTXCLKTOPLBUFG(),
        .FMIOGEM0SIGNALDETECT(),
        .FMIOGEM1FIFORXCLKFROMPL(),
        .FMIOGEM1FIFORXCLKTOPLBUFG(),
        .FMIOGEM1FIFOTXCLKFROMPL(),
        .FMIOGEM1FIFOTXCLKTOPLBUFG(),
        .FMIOGEM1SIGNALDETECT(),
        .FMIOGEM2FIFORXCLKFROMPL(),
        .FMIOGEM2FIFORXCLKTOPLBUFG(),
        .FMIOGEM2FIFOTXCLKFROMPL(),
        .FMIOGEM2FIFOTXCLKTOPLBUFG(),
        .FMIOGEM2SIGNALDETECT(),
        .FMIOGEM3FIFORXCLKFROMPL(),
        .FMIOGEM3FIFORXCLKTOPLBUFG(),
        .FMIOGEM3FIFOTXCLKFROMPL(),
        .FMIOGEM3FIFOTXCLKTOPLBUFG(),
        .FMIOGEM3SIGNALDETECT(),
        .FMIOGEMTSUCLKFROMPL(),
        .FMIOGEMTSUCLKTOPLBUFG(),
        .FTMGPI(),
        .FTMGPO(),
        .GDMA2PLCACK(),
        .GDMA2PLTVLD(),
        .GDMAFCICLK(),
        .MAXIGP0ACLK(),
        .MAXIGP0ARADDR(),
        .MAXIGP0ARBURST(),
        .MAXIGP0ARCACHE(),
        .MAXIGP0ARID(),
        .MAXIGP0ARLEN(),
        .MAXIGP0ARLOCK(),
        .MAXIGP0ARPROT(),
        .MAXIGP0ARQOS(),
        .MAXIGP0ARREADY(),
        .MAXIGP0ARSIZE(),
        .MAXIGP0ARUSER(),
        .MAXIGP0ARVALID(),
        .MAXIGP0AWADDR(),
        .MAXIGP0AWBURST(),
        .MAXIGP0AWCACHE(),
        .MAXIGP0AWID(),
        .MAXIGP0AWLEN(),
        .MAXIGP0AWLOCK(),
        .MAXIGP0AWPROT(),
        .MAXIGP0AWQOS(),
        .MAXIGP0AWREADY(),
        .MAXIGP0AWSIZE(),
        .MAXIGP0AWUSER(),
        .MAXIGP0AWVALID(),
        .MAXIGP0BID(),
        .MAXIGP0BREADY(),
        .MAXIGP0BRESP(),
        .MAXIGP0BVALID(),
        .MAXIGP0RDATA(),
        .MAXIGP0RID(),
        .MAXIGP0RLAST(),
        .MAXIGP0RREADY(),
        .MAXIGP0RRESP(),
        .MAXIGP0RVALID(),
        .MAXIGP0WDATA(),
        .MAXIGP0WLAST(),
        .MAXIGP0WREADY(),
        .MAXIGP0WSTRB(),
        .MAXIGP0WVALID(),
        .MAXIGP1ACLK(),
        .MAXIGP1ARADDR(),
        .MAXIGP1ARBURST(),
        .MAXIGP1ARCACHE(),
        .MAXIGP1ARID(),
        .MAXIGP1ARLEN(),
        .MAXIGP1ARLOCK(),
        .MAXIGP1ARPROT(),
        .MAXIGP1ARQOS(),
        .MAXIGP1ARREADY(),
        .MAXIGP1ARSIZE(),
        .MAXIGP1ARUSER(),
        .MAXIGP1ARVALID(),
        .MAXIGP1AWADDR(),
        .MAXIGP1AWBURST(),
        .MAXIGP1AWCACHE(),
        .MAXIGP1AWID(),
        .MAXIGP1AWLEN(),
        .MAXIGP1AWLOCK(),
        .MAXIGP1AWPROT(),
        .MAXIGP1AWQOS(),
        .MAXIGP1AWREADY(),
        .MAXIGP1AWSIZE(),
        .MAXIGP1AWUSER(),
        .MAXIGP1AWVALID(),
        .MAXIGP1BID(),
        .MAXIGP1BREADY(),
        .MAXIGP1BRESP(),
        .MAXIGP1BVALID(),
        .MAXIGP1RDATA(),
        .MAXIGP1RID(),
        .MAXIGP1RLAST(),
        .MAXIGP1RREADY(),
        .MAXIGP1RRESP(),
        .MAXIGP1RVALID(),
        .MAXIGP1WDATA(),
        .MAXIGP1WLAST(),
        .MAXIGP1WREADY(),
        .MAXIGP1WSTRB(),
        .MAXIGP1WVALID(),
        .MAXIGP2ACLK(),
        .MAXIGP2ARADDR(),
        .MAXIGP2ARBURST(),
        .MAXIGP2ARCACHE(),
        .MAXIGP2ARID(),
        .MAXIGP2ARLEN(),
        .MAXIGP2ARLOCK(),
        .MAXIGP2ARPROT(),
        .MAXIGP2ARQOS(),
        .MAXIGP2ARREADY(),
        .MAXIGP2ARSIZE(),
        .MAXIGP2ARUSER(),
        .MAXIGP2ARVALID(),
        .MAXIGP2AWADDR(),
        .MAXIGP2AWBURST(),
        .MAXIGP2AWCACHE(),
        .MAXIGP2AWID(),
        .MAXIGP2AWLEN(),
        .MAXIGP2AWLOCK(),
        .MAXIGP2AWPROT(),
        .MAXIGP2AWQOS(),
        .MAXIGP2AWREADY(),
        .MAXIGP2AWSIZE(),
        .MAXIGP2AWUSER(),
        .MAXIGP2AWVALID(),
        .MAXIGP2BID(),
        .MAXIGP2BREADY(),
        .MAXIGP2BRESP(),
        .MAXIGP2BVALID(),
        .MAXIGP2RDATA(),
        .MAXIGP2RID(),
        .MAXIGP2RLAST(),
        .MAXIGP2RREADY(),
        .MAXIGP2RRESP(),
        .MAXIGP2RVALID(),
        .MAXIGP2WDATA(),
        .MAXIGP2WLAST(),
        .MAXIGP2WREADY(),
        .MAXIGP2WSTRB(),
        .MAXIGP2WVALID(),
        .NFIQ0LPDRPU(),
        .NFIQ1LPDRPU(),
        .NIRQ0LPDRPU(),
        .NIRQ1LPDRPU(),
        .OSCRTCCLK(),
        .PL2ADMACVLD(),
        .PL2ADMATACK(),
        .PL2GDMACVLD(),
        .PL2GDMATACK(),
        .PLACECLK(),
        .PLACPINACT(),
        .PLCLK({pl_clk3,pl_clk2,pl_clk1,pl_clk_unbuffered}),
        .PLFPGASTOP(),
        .PLLAUXREFCLKFPD(),
        .PLLAUXREFCLKLPD(),
        .PLPMUGPI(),
        .PLPSAPUGICFIQ(),
        .PLPSAPUGICIRQ(),
        .PLPSEVENTI(),
        .PLPSIRQ0(),
        .PLPSIRQ1(),
        .PLPSTRACECLK(),
        .PLPSTRIGACK(),
        .PLPSTRIGGER(),
        .PMUAIBAFIFMFPDREQ(),
        .PMUAIBAFIFMLPDREQ(),
        .PMUERRORFROMPL(),
        .PMUERRORTOPL(),
        .PMUPLGPO(),
        .PSPLEVENTO(),
        .PSPLIRQFPD(),
        .PSPLIRQLPD(),
        .PSPLSTANDBYWFE(),
        .PSPLSTANDBYWFI(),
        .PSPLTRACECTL(),
        .PSPLTRACEDATA(),
        .PSPLTRIGACK(),
        .PSPLTRIGGER(),
        .PSS_ALTO_CORE_PAD_BOOTMODE(),
        .PSS_ALTO_CORE_PAD_CLK(),
        .PSS_ALTO_CORE_PAD_DONEB(),
        .PSS_ALTO_CORE_PAD_DRAMA(),
        .PSS_ALTO_CORE_PAD_DRAMACTN(),
        .PSS_ALTO_CORE_PAD_DRAMALERTN(),
        .PSS_ALTO_CORE_PAD_DRAMBA(),
        .PSS_ALTO_CORE_PAD_DRAMBG(),
        .PSS_ALTO_CORE_PAD_DRAMCK(),
        .PSS_ALTO_CORE_PAD_DRAMCKE(),
        .PSS_ALTO_CORE_PAD_DRAMCKN(),
        .PSS_ALTO_CORE_PAD_DRAMCSN(),
        .PSS_ALTO_CORE_PAD_DRAMDM(),
        .PSS_ALTO_CORE_PAD_DRAMDQ(),
        .PSS_ALTO_CORE_PAD_DRAMDQS(),
        .PSS_ALTO_CORE_PAD_DRAMDQSN(),
        .PSS_ALTO_CORE_PAD_DRAMODT(),
        .PSS_ALTO_CORE_PAD_DRAMPARITY(),
        .PSS_ALTO_CORE_PAD_DRAMRAMRSTN(),
        .PSS_ALTO_CORE_PAD_ERROROUT(),
        .PSS_ALTO_CORE_PAD_ERRORSTATUS(),
        .PSS_ALTO_CORE_PAD_INITB(),
        .PSS_ALTO_CORE_PAD_JTAGTCK(),
        .PSS_ALTO_CORE_PAD_JTAGTDI(),
        .PSS_ALTO_CORE_PAD_JTAGTDO(),
        .PSS_ALTO_CORE_PAD_JTAGTMS(),
        .PSS_ALTO_CORE_PAD_MGTRXN0IN(),
        .PSS_ALTO_CORE_PAD_MGTRXN1IN(),
        .PSS_ALTO_CORE_PAD_MGTRXN2IN(),
        .PSS_ALTO_CORE_PAD_MGTRXN3IN(),
        .PSS_ALTO_CORE_PAD_MGTRXP0IN(),
        .PSS_ALTO_CORE_PAD_MGTRXP1IN(),
        .PSS_ALTO_CORE_PAD_MGTRXP2IN(),
        .PSS_ALTO_CORE_PAD_MGTRXP3IN(),
        .PSS_ALTO_CORE_PAD_MGTTXN0OUT(),
        .PSS_ALTO_CORE_PAD_MGTTXN1OUT(),
        .PSS_ALTO_CORE_PAD_MGTTXN2OUT(),
        .PSS_ALTO_CORE_PAD_MGTTXN3OUT(),
        .PSS_ALTO_CORE_PAD_MGTTXP0OUT(),
        .PSS_ALTO_CORE_PAD_MGTTXP1OUT(),
        .PSS_ALTO_CORE_PAD_MGTTXP2OUT(),
        .PSS_ALTO_CORE_PAD_MGTTXP3OUT(),
        .PSS_ALTO_CORE_PAD_MIO(),
        .PSS_ALTO_CORE_PAD_PADI(),
        .PSS_ALTO_CORE_PAD_PADO(),
        .PSS_ALTO_CORE_PAD_PORB(),
        .PSS_ALTO_CORE_PAD_PROGB(),
        .PSS_ALTO_CORE_PAD_RCALIBINOUT(),
        .PSS_ALTO_CORE_PAD_REFN0IN(),
        .PSS_ALTO_CORE_PAD_REFN1IN(),
        .PSS_ALTO_CORE_PAD_REFN2IN(),
        .PSS_ALTO_CORE_PAD_REFN3IN(),
        .PSS_ALTO_CORE_PAD_REFP0IN(),
        .PSS_ALTO_CORE_PAD_REFP1IN(),
        .PSS_ALTO_CORE_PAD_REFP2IN(),
        .PSS_ALTO_CORE_PAD_REFP3IN(),
        .PSS_ALTO_CORE_PAD_SRSTB(),
        .PSS_ALTO_CORE_PAD_ZQ(),
        .RPUEVENTI0(),
        .RPUEVENTI1(),
        .RPUEVENTO0(),
        .RPUEVENTO1(),
        .SACEFPDACADDR(),
        .SACEFPDACPROT(),
        .SACEFPDACREADY(),
        .SACEFPDACSNOOP(),
        .SACEFPDACVALID(),
        .SACEFPDARADDR(),
        .SACEFPDARBAR(),
        .SACEFPDARBURST(),
        .SACEFPDARCACHE(),
        .SACEFPDARDOMAIN(),
        .SACEFPDARID(),
        .SACEFPDARLEN(),
        .SACEFPDARLOCK(),
        .SACEFPDARPROT(),
        .SACEFPDARQOS(),
        .SACEFPDARREADY(),
        .SACEFPDARREGION(),
        .SACEFPDARSIZE(),
        .SACEFPDARSNOOP(),
        .SACEFPDARUSER(),
        .SACEFPDARVALID(),
        .SACEFPDAWADDR(),
        .SACEFPDAWBAR(),
        .SACEFPDAWBURST(),
        .SACEFPDAWCACHE(),
        .SACEFPDAWDOMAIN(),
        .SACEFPDAWID(),
        .SACEFPDAWLEN(),
        .SACEFPDAWLOCK(),
        .SACEFPDAWPROT(),
        .SACEFPDAWQOS(),
        .SACEFPDAWREADY(),
        .SACEFPDAWREGION(),
        .SACEFPDAWSIZE(),
        .SACEFPDAWSNOOP(),
        .SACEFPDAWUSER(),
        .SACEFPDAWVALID(),
        .SACEFPDBID(),
        .SACEFPDBREADY(),
        .SACEFPDBRESP(),
        .SACEFPDBUSER(),
        .SACEFPDBVALID(),
        .SACEFPDCDDATA(),
        .SACEFPDCDLAST(),
        .SACEFPDCDREADY(),
        .SACEFPDCDVALID(),
        .SACEFPDCRREADY(),
        .SACEFPDCRRESP(),
        .SACEFPDCRVALID(),
        .SACEFPDRACK(),
        .SACEFPDRDATA(),
        .SACEFPDRID(),
        .SACEFPDRLAST(),
        .SACEFPDRREADY(),
        .SACEFPDRRESP(),
        .SACEFPDRUSER(),
        .SACEFPDRVALID(),
        .SACEFPDWACK(),
        .SACEFPDWDATA(),
        .SACEFPDWLAST(),
        .SACEFPDWREADY(),
        .SACEFPDWSTRB(),
        .SACEFPDWUSER(),
        .SACEFPDWVALID(),
        .SAXIACPACLK(),
        .SAXIACPARADDR(),
        .SAXIACPARBURST(),
        .SAXIACPARCACHE(),
        .SAXIACPARID(),
        .SAXIACPARLEN(),
        .SAXIACPARLOCK(),
        .SAXIACPARPROT(),
        .SAXIACPARQOS(),
        .SAXIACPARREADY(),
        .SAXIACPARSIZE(),
        .SAXIACPARUSER(),
        .SAXIACPARVALID(),
        .SAXIACPAWADDR(),
        .SAXIACPAWBURST(),
        .SAXIACPAWCACHE(),
        .SAXIACPAWID(),
        .SAXIACPAWLEN(),
        .SAXIACPAWLOCK(),
        .SAXIACPAWPROT(),
        .SAXIACPAWQOS(),
        .SAXIACPAWREADY(),
        .SAXIACPAWSIZE(),
        .SAXIACPAWUSER(),
        .SAXIACPAWVALID(),
        .SAXIACPBID(),
        .SAXIACPBREADY(),
        .SAXIACPBRESP(),
        .SAXIACPBVALID(),
        .SAXIACPRDATA(),
        .SAXIACPRID(),
        .SAXIACPRLAST(),
        .SAXIACPRREADY(),
        .SAXIACPRRESP(),
        .SAXIACPRVALID(),
        .SAXIACPWDATA(),
        .SAXIACPWLAST(),
        .SAXIACPWREADY(),
        .SAXIACPWSTRB(),
        .SAXIACPWVALID(),
        .SAXIGP0ARADDR(),
        .SAXIGP0ARBURST(),
        .SAXIGP0ARCACHE(),
        .SAXIGP0ARID(),
        .SAXIGP0ARLEN(),
        .SAXIGP0ARLOCK(),
        .SAXIGP0ARPROT(),
        .SAXIGP0ARQOS(),
        .SAXIGP0ARREADY(),
        .SAXIGP0ARSIZE(),
        .SAXIGP0ARUSER(),
        .SAXIGP0ARVALID(),
        .SAXIGP0AWADDR(),
        .SAXIGP0AWBURST(),
        .SAXIGP0AWCACHE(),
        .SAXIGP0AWID(),
        .SAXIGP0AWLEN(),
        .SAXIGP0AWLOCK(),
        .SAXIGP0AWPROT(),
        .SAXIGP0AWQOS(),
        .SAXIGP0AWREADY(),
        .SAXIGP0AWSIZE(),
        .SAXIGP0AWUSER(),
        .SAXIGP0AWVALID(),
        .SAXIGP0BID(),
        .SAXIGP0BREADY(),
        .SAXIGP0BRESP(),
        .SAXIGP0BVALID(),
        .SAXIGP0RACOUNT(),
        .SAXIGP0RCLK(),
        .SAXIGP0RCOUNT(),
        .SAXIGP0RDATA(),
        .SAXIGP0RID(),
        .SAXIGP0RLAST(),
        .SAXIGP0RREADY(),
        .SAXIGP0RRESP(),
        .SAXIGP0RVALID(),
        .SAXIGP0WACOUNT(),
        .SAXIGP0WCLK(),
        .SAXIGP0WCOUNT(),
        .SAXIGP0WDATA(),
        .SAXIGP0WLAST(),
        .SAXIGP0WREADY(),
        .SAXIGP0WSTRB(),
        .SAXIGP0WVALID(),
        .SAXIGP1ARADDR(),
        .SAXIGP1ARBURST(),
        .SAXIGP1ARCACHE(),
        .SAXIGP1ARID(),
        .SAXIGP1ARLEN(),
        .SAXIGP1ARLOCK(),
        .SAXIGP1ARPROT(),
        .SAXIGP1ARQOS(),
        .SAXIGP1ARREADY(),
        .SAXIGP1ARSIZE(),
        .SAXIGP1ARUSER(),
        .SAXIGP1ARVALID(),
        .SAXIGP1AWADDR(),
        .SAXIGP1AWBURST(),
        .SAXIGP1AWCACHE(),
        .SAXIGP1AWID(),
        .SAXIGP1AWLEN(),
        .SAXIGP1AWLOCK(),
        .SAXIGP1AWPROT(),
        .SAXIGP1AWQOS(),
        .SAXIGP1AWREADY(),
        .SAXIGP1AWSIZE(),
        .SAXIGP1AWUSER(),
        .SAXIGP1AWVALID(),
        .SAXIGP1BID(),
        .SAXIGP1BREADY(),
        .SAXIGP1BRESP(),
        .SAXIGP1BVALID(),
        .SAXIGP1RACOUNT(),
        .SAXIGP1RCLK(),
        .SAXIGP1RCOUNT(),
        .SAXIGP1RDATA(),
        .SAXIGP1RID(),
        .SAXIGP1RLAST(),
        .SAXIGP1RREADY(),
        .SAXIGP1RRESP(),
        .SAXIGP1RVALID(),
        .SAXIGP1WACOUNT(),
        .SAXIGP1WCLK(),
        .SAXIGP1WCOUNT(),
        .SAXIGP1WDATA(),
        .SAXIGP1WLAST(),
        .SAXIGP1WREADY(),
        .SAXIGP1WSTRB(),
        .SAXIGP1WVALID(),
        .SAXIGP2ARADDR(),
        .SAXIGP2ARBURST(),
        .SAXIGP2ARCACHE(),
        .SAXIGP2ARID(),
        .SAXIGP2ARLEN(),
        .SAXIGP2ARLOCK(),
        .SAXIGP2ARPROT(),
        .SAXIGP2ARQOS(),
        .SAXIGP2ARREADY(),
        .SAXIGP2ARSIZE(),
        .SAXIGP2ARUSER(),
        .SAXIGP2ARVALID(),
        .SAXIGP2AWADDR(),
        .SAXIGP2AWBURST(),
        .SAXIGP2AWCACHE(),
        .SAXIGP2AWID(),
        .SAXIGP2AWLEN(),
        .SAXIGP2AWLOCK(),
        .SAXIGP2AWPROT(),
        .SAXIGP2AWQOS(),
        .SAXIGP2AWREADY(),
        .SAXIGP2AWSIZE(),
        .SAXIGP2AWUSER(),
        .SAXIGP2AWVALID(),
        .SAXIGP2BID(),
        .SAXIGP2BREADY(),
        .SAXIGP2BRESP(),
        .SAXIGP2BVALID(),
        .SAXIGP2RACOUNT(),
        .SAXIGP2RCLK(),
        .SAXIGP2RCOUNT(),
        .SAXIGP2RDATA(),
        .SAXIGP2RID(),
        .SAXIGP2RLAST(),
        .SAXIGP2RREADY(),
        .SAXIGP2RRESP(),
        .SAXIGP2RVALID(),
        .SAXIGP2WACOUNT(),
        .SAXIGP2WCLK(),
        .SAXIGP2WCOUNT(),
        .SAXIGP2WDATA(),
        .SAXIGP2WLAST(),
        .SAXIGP2WREADY(),
        .SAXIGP2WSTRB(),
        .SAXIGP2WVALID(),
        .SAXIGP3ARADDR(),
        .SAXIGP3ARBURST(),
        .SAXIGP3ARCACHE(),
        .SAXIGP3ARID(),
        .SAXIGP3ARLEN(),
        .SAXIGP3ARLOCK(),
        .SAXIGP3ARPROT(),
        .SAXIGP3ARQOS(),
        .SAXIGP3ARREADY(),
        .SAXIGP3ARSIZE(),
        .SAXIGP3ARUSER(),
        .SAXIGP3ARVALID(),
        .SAXIGP3AWADDR(),
        .SAXIGP3AWBURST(),
        .SAXIGP3AWCACHE(),
        .SAXIGP3AWID(),
        .SAXIGP3AWLEN(),
        .SAXIGP3AWLOCK(),
        .SAXIGP3AWPROT(),
        .SAXIGP3AWQOS(),
        .SAXIGP3AWREADY(),
        .SAXIGP3AWSIZE(),
        .SAXIGP3AWUSER(),
        .SAXIGP3AWVALID(),
        .SAXIGP3BID(),
        .SAXIGP3BREADY(),
        .SAXIGP3BRESP(),
        .SAXIGP3BVALID(),
        .SAXIGP3RACOUNT(),
        .SAXIGP3RCLK(),
        .SAXIGP3RCOUNT(),
        .SAXIGP3RDATA(),
        .SAXIGP3RID(),
        .SAXIGP3RLAST(),
        .SAXIGP3RREADY(),
        .SAXIGP3RRESP(),
        .SAXIGP3RVALID(),
        .SAXIGP3WACOUNT(),
        .SAXIGP3WCLK(),
        .SAXIGP3WCOUNT(),
        .SAXIGP3WDATA(),
        .SAXIGP3WLAST(),
        .SAXIGP3WREADY(),
        .SAXIGP3WSTRB(),
        .SAXIGP3WVALID(),
        .SAXIGP4ARADDR(),
        .SAXIGP4ARBURST(),
        .SAXIGP4ARCACHE(),
        .SAXIGP4ARID(),
        .SAXIGP4ARLEN(),
        .SAXIGP4ARLOCK(),
        .SAXIGP4ARPROT(),
        .SAXIGP4ARQOS(),
        .SAXIGP4ARREADY(),
        .SAXIGP4ARSIZE(),
        .SAXIGP4ARUSER(),
        .SAXIGP4ARVALID(),
        .SAXIGP4AWADDR(),
        .SAXIGP4AWBURST(),
        .SAXIGP4AWCACHE(),
        .SAXIGP4AWID(),
        .SAXIGP4AWLEN(),
        .SAXIGP4AWLOCK(),
        .SAXIGP4AWPROT(),
        .SAXIGP4AWQOS(),
        .SAXIGP4AWREADY(),
        .SAXIGP4AWSIZE(),
        .SAXIGP4AWUSER(),
        .SAXIGP4AWVALID(),
        .SAXIGP4BID(),
        .SAXIGP4BREADY(),
        .SAXIGP4BRESP(),
        .SAXIGP4BVALID(),
        .SAXIGP4RACOUNT(),
        .SAXIGP4RCLK(),
        .SAXIGP4RCOUNT(),
        .SAXIGP4RDATA(),
        .SAXIGP4RID(),
        .SAXIGP4RLAST(),
        .SAXIGP4RREADY(),
        .SAXIGP4RRESP(),
        .SAXIGP4RVALID(),
        .SAXIGP4WACOUNT(),
        .SAXIGP4WCLK(),
        .SAXIGP4WCOUNT(),
        .SAXIGP4WDATA(),
        .SAXIGP4WLAST(),
        .SAXIGP4WREADY(),
        .SAXIGP4WSTRB(),
        .SAXIGP4WVALID(),
        .SAXIGP5ARADDR(),
        .SAXIGP5ARBURST(),
        .SAXIGP5ARCACHE(),
        .SAXIGP5ARID(),
        .SAXIGP5ARLEN(),
        .SAXIGP5ARLOCK(),
        .SAXIGP5ARPROT(),
        .SAXIGP5ARQOS(),
        .SAXIGP5ARREADY(),
        .SAXIGP5ARSIZE(),
        .SAXIGP5ARUSER(),
        .SAXIGP5ARVALID(),
        .SAXIGP5AWADDR(),
        .SAXIGP5AWBURST(),
        .SAXIGP5AWCACHE(),
        .SAXIGP5AWID(),
        .SAXIGP5AWLEN(),
        .SAXIGP5AWLOCK(),
        .SAXIGP5AWPROT(),
        .SAXIGP5AWQOS(),
        .SAXIGP5AWREADY(),
        .SAXIGP5AWSIZE(),
        .SAXIGP5AWUSER(),
        .SAXIGP5AWVALID(),
        .SAXIGP5BID(),
        .SAXIGP5BREADY(),
        .SAXIGP5BRESP(),
        .SAXIGP5BVALID(),
        .SAXIGP5RACOUNT(),
        .SAXIGP5RCLK(),
        .SAXIGP5RCOUNT(),
        .SAXIGP5RDATA(),
        .SAXIGP5RID(),
        .SAXIGP5RLAST(),
        .SAXIGP5RREADY(),
        .SAXIGP5RRESP(),
        .SAXIGP5RVALID(),
        .SAXIGP5WACOUNT(),
        .SAXIGP5WCLK(),
        .SAXIGP5WCOUNT(),
        .SAXIGP5WDATA(),
        .SAXIGP5WLAST(),
        .SAXIGP5WREADY(),
        .SAXIGP5WSTRB(),
        .SAXIGP5WVALID(),
        .SAXIGP6ARADDR(),
        .SAXIGP6ARBURST(),
        .SAXIGP6ARCACHE(),
        .SAXIGP6ARID(),
        .SAXIGP6ARLEN(),
        .SAXIGP6ARLOCK(),
        .SAXIGP6ARPROT(),
        .SAXIGP6ARQOS(),
        .SAXIGP6ARREADY(),
        .SAXIGP6ARSIZE(),
        .SAXIGP6ARUSER(),
        .SAXIGP6ARVALID(),
        .SAXIGP6AWADDR(),
        .SAXIGP6AWBURST(),
        .SAXIGP6AWCACHE(),
        .SAXIGP6AWID(),
        .SAXIGP6AWLEN(),
        .SAXIGP6AWLOCK(),
        .SAXIGP6AWPROT(),
        .SAXIGP6AWQOS(),
        .SAXIGP6AWREADY(),
        .SAXIGP6AWSIZE(),
        .SAXIGP6AWUSER(),
        .SAXIGP6AWVALID(),
        .SAXIGP6BID(),
        .SAXIGP6BREADY(),
        .SAXIGP6BRESP(),
        .SAXIGP6BVALID(),
        .SAXIGP6RACOUNT(),
        .SAXIGP6RCLK(),
        .SAXIGP6RCOUNT(),
        .SAXIGP6RDATA(),
        .SAXIGP6RID(),
        .SAXIGP6RLAST(),
        .SAXIGP6RREADY(),
        .SAXIGP6RRESP(),
        .SAXIGP6RVALID(),
        .SAXIGP6WACOUNT(),
        .SAXIGP6WCLK(),
        .SAXIGP6WCOUNT(),
        .SAXIGP6WDATA(),
        .SAXIGP6WLAST(),
        .SAXIGP6WREADY(),
        .SAXIGP6WSTRB(),
        .SAXIGP6WVALID(),
        .STMEVENT());
  VCC VCC
       (.P(\<const1> ));
  (* BOX_TYPE = "PRIMITIVE" *)
  BUFG_PS #(
    .SIM_DEVICE("ULTRASCALE_PLUS"),
    .STARTUP_SYNC("FALSE"))
    \buffer_pl_clk_0.PL_CLK_0_BUFG
       (.I(pl_clk_unbuffered),
        .O(pl_clk0));


endmodule
